`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:40:07 01/29/2022 
// Design Name: 
// Module Name:    keypad4x4 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module keypad4x4(
    input clk,
    input [3:0] row,
    output [3:0] col,
    output [3:0] hex,
    output keydown
    );


endmodule
